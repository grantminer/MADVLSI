* NGSPICE file created from bias.ext - technology: sky130A

X0 Vcp Ib Vbp Vcp sky130_fd_pr__nfet_01v8 ad=6 pd=25 as=3 ps=12.5 w=12 l=0.5
X1 a_700_0# Ib a_500_0# Vcp sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X2 a_n100_8040# a_n100_8040# a_100_5330# Vcp sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X3 a_2450_8040# Vbp Vcn Vcn sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X4 a_n100_8040# a_n100_8040# a_100_5330# Vcp sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X5 a_1000_5300# a_1000_5300# a_100_5330# Vcp sky130_fd_pr__nfet_01v8 ad=6 pd=25 as=3 ps=12.5 w=12 l=0.5
X6 Vcp Ib a_n100_0# Vcp sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=6 ps=25 w=12 l=0.5
X7 a_2850_8040# Vbp a_2650_8040# Vcn sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X8 a_200_2600# a_200_2600# a_100_2660# Vcn sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X9 a_200_2600# a_200_2600# a_100_2660# Vcn sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X10 Vcn a_200_2600# a_100_2660# Vcn sky130_fd_pr__pfet_01v8 ad=6 pd=25 as=3 ps=12.5 w=12 l=0.5
X11 Vcp a_2350_5300# a_2250_5330# Vcp sky130_fd_pr__nfet_01v8 ad=6 pd=25 as=3 ps=12.5 w=12 l=0.5
X12 a_2250_0# Ib a_2050_0# Vcp sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=6 ps=25 w=12 l=0.5
X13 Vcp Ib Ib Vcp sky130_fd_pr__nfet_01v8 ad=6 pd=25 as=3 ps=12.5 w=12 l=0.5
X14 a_2850_0# Ib a_2650_0# Vcp sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X15 a_2250_5330# a_2050_5330# a_2050_5330# Vcp sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=6 ps=25 w=12 l=0.5
X16 a_3150_2600# a_3150_2600# a_2250_2660# Vcn sky130_fd_pr__pfet_01v8 ad=6 pd=25 as=3 ps=12.5 w=12 l=0.5
X17 a_2250_5330# a_2350_5300# a_2350_5300# Vcp sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X18 a_2250_5330# a_2350_5300# a_2350_5300# Vcp sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X19 a_2250_2660# a_2050_0# Vcn Vcn sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=6 ps=25 w=12 l=0.5
X20 a_300_0# Ib Vcp Vcp sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X21 Vbp Vbp Vcn Vcn sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=6 ps=25 w=12 l=0.5
X22 a_2250_2660# a_2050_0# a_2050_0# Vcn sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X23 a_300_8040# Vbp a_100_8040# Vcn sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X24 a_2250_2660# a_2050_0# a_2050_0# Vcn sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X25 a_900_0# Ib a_700_0# Vcp sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X26 a_700_8040# Vbp a_500_8040# Vcn sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X27 a_1000_5300# Vbp Vcn Vcn sky130_fd_pr__pfet_01v8 ad=6 pd=25 as=3 ps=12.5 w=12 l=0.5
X28 a_200_2600# Ib a_900_0# Vcp sky130_fd_pr__nfet_01v8 ad=6 pd=25 as=3 ps=12.5 w=12 l=0.5
X29 Vbp Ib Vcp Vcp sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=6 ps=25 w=12 l=0.5
X30 a_2350_5300# Vbp a_3050_8040# Vcn sky130_fd_pr__pfet_01v8 ad=6 pd=25 as=3 ps=12.5 w=12 l=0.5
X31 a_2450_0# Ib a_2250_0# Vcp sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X32 a_100_5330# a_n100_8040# Vcp Vcp sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=6 ps=25 w=12 l=0.5
X33 a_100_5330# a_n100_8040# a_n100_8040# Vcp sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X34 Vcp Ib a_2850_0# Vcp sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X35 Vcn Vbp a_2050_5330# Vcn sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=6 ps=25 w=12 l=0.5
X36 a_2650_8040# Vbp a_2450_8040# Vcn sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X37 a_100_5330# a_n100_8040# a_n100_8040# Vcp sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X38 a_3050_8040# Vbp a_2850_8040# Vcn sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X39 a_100_2660# a_n100_0# a_n100_0# Vcn sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=6 ps=25 w=12 l=0.5
X40 a_100_2660# a_200_2600# a_200_2600# Vcn sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X41 a_100_2660# a_200_2600# a_200_2600# Vcn sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X42 a_500_0# Ib a_300_0# Vcp sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X43 a_2350_5300# a_2350_5300# a_2250_5330# Vcp sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X44 a_2350_5300# a_2350_5300# a_2250_5330# Vcp sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X45 Vcn Vbp Vbp Vcn sky130_fd_pr__pfet_01v8 ad=6 pd=25 as=3 ps=12.5 w=12 l=0.5
X46 a_2050_0# a_2050_0# a_2250_2660# Vcn sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X47 a_2050_0# a_2050_0# a_2250_2660# Vcn sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X48 Ib Ib Vcp Vcp sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=6 ps=25 w=12 l=0.5
X49 a_2650_0# Ib a_2450_0# Vcp sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X50 a_100_8040# Vbp a_n100_8040# Vcn sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=6 ps=25 w=12 l=0.5
X51 a_500_8040# Vbp a_300_8040# Vcn sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X52 Vcn Vbp a_700_8040# Vcn sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X53 a_3150_2600# Ib Vcp Vcp sky130_fd_pr__nfet_01v8 ad=6 pd=25 as=3 ps=12.5 w=12 l=0.5

