magic
tech sky130A
timestamp 1697738063
<< poly >>
rect 265 7385 315 7395
rect 265 7355 275 7385
rect 305 7355 315 7385
rect 265 7345 315 7355
rect 265 6000 315 6010
rect 265 5970 275 6000
rect 305 5970 315 6000
rect 265 5960 315 5970
rect -40 5690 10 5700
rect -40 5660 -30 5690
rect 0 5660 10 5690
rect -40 5545 10 5660
rect -40 5515 -30 5545
rect 0 5515 10 5545
rect -40 5505 10 5515
rect -235 5415 150 5425
rect -235 5385 110 5415
rect 140 5385 150 5415
rect -235 5375 150 5385
rect 265 4665 315 4675
rect 265 4635 275 4665
rect 305 4635 315 4665
rect 265 4625 315 4635
rect 245 2650 320 2660
rect 245 2620 255 2650
rect 285 2645 320 2650
rect 285 2620 295 2645
rect 245 2610 295 2620
rect -120 1395 220 1405
rect -120 1390 180 1395
rect -185 1365 180 1390
rect 210 1365 220 1395
rect -185 1355 220 1365
rect 265 1235 315 1245
rect 265 1205 275 1235
rect 305 1205 315 1235
rect 265 1195 315 1205
rect -40 -100 150 -90
rect -40 -130 -30 -100
rect 0 -130 110 -100
rect 140 -130 150 -100
rect -40 -140 150 -130
rect 265 -100 315 -90
rect 265 -130 275 -100
rect 305 -130 315 -100
rect 265 -140 315 -130
rect 265 -1510 315 -1500
rect 265 -1540 275 -1510
rect 305 -1540 315 -1510
rect 265 -1550 315 -1540
<< polycont >>
rect 275 7355 305 7385
rect 275 5970 305 6000
rect -30 5660 0 5690
rect -30 5515 0 5545
rect 110 5385 140 5415
rect 275 4635 305 4665
rect 255 2620 285 2650
rect 180 1365 210 1395
rect 275 1205 305 1235
rect -30 -130 0 -100
rect 110 -130 140 -100
rect 275 -130 305 -100
rect 275 -1540 305 -1510
<< locali >>
rect -780 7385 315 7395
rect -780 7355 275 7385
rect 305 7355 315 7385
rect -780 7345 315 7355
rect -780 5625 -740 7345
rect -40 6000 315 6010
rect -40 5970 275 6000
rect 305 5970 315 6000
rect -40 5960 315 5970
rect -40 5690 10 5960
rect -40 5660 -30 5690
rect 0 5660 10 5690
rect -40 5650 10 5660
rect -785 5575 80 5625
rect -780 5460 -740 5575
rect -40 5545 10 5555
rect -40 5515 -30 5545
rect 0 5515 10 5545
rect -40 1400 10 5515
rect -55 1380 10 1400
rect -1020 40 -980 70
rect -1940 -10 -980 40
rect -40 -100 10 1380
rect -40 -130 -30 -100
rect 0 -130 10 -100
rect -40 -140 10 -130
rect 30 -1500 80 5575
rect 100 5415 150 5425
rect 100 5385 110 5415
rect 140 5385 150 5415
rect 100 4675 150 5385
rect 100 4665 315 4675
rect 100 4635 275 4665
rect 305 4635 315 4665
rect 100 4625 315 4635
rect 100 1245 150 4625
rect 170 2650 295 2660
rect 170 2620 255 2650
rect 285 2620 295 2650
rect 170 2610 295 2620
rect 170 1395 220 2610
rect 170 1365 180 1395
rect 210 1365 220 1395
rect 170 1355 220 1365
rect 100 1235 315 1245
rect 100 1205 275 1235
rect 305 1205 315 1235
rect 100 1195 315 1205
rect 825 1140 1000 1160
rect 100 -100 315 -90
rect 100 -130 110 -100
rect 140 -130 275 -100
rect 305 -130 315 -100
rect 100 -140 315 -130
rect 30 -1510 315 -1500
rect 30 -1540 275 -1510
rect 305 -1540 315 -1510
rect 30 -1550 315 -1540
<< metal1 >>
rect -1880 7395 880 7465
rect -1880 5455 385 7395
rect 840 7380 880 7395
rect -185 1355 -55 1395
rect -1940 -1550 425 60
use bias  bias_0
timestamp 1697565880
transform 1 0 -1810 0 1 140
box -130 -80 1755 5320
use fcda  fcda_0
timestamp 1697505651
transform 1 0 539 0 1 -2289
box -224 739 457 9684
<< labels >>
rlabel locali -1940 15 -1940 15 7 Ib
port 1 w
rlabel locali 1000 1150 1000 1150 3 Vout
port 2 e
rlabel metal1 -385 7465 -385 7465 1 VP
port 3 n
rlabel metal1 -570 -1550 -570 -1550 5 VN
port 4 s
<< end >>
