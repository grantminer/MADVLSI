magic
tech sky130A
magscale 1 2
timestamp 1695946031
<< nwell >>
rect -226 946 556 1978
<< nmos >>
rect -90 60 -60 862
rect 62 662 92 862
rect 214 662 244 862
rect 366 662 396 862
rect 62 60 92 260
rect 214 60 244 260
rect 346 60 376 260
<< pmos >>
rect -90 1584 -60 1784
rect 42 1584 72 1784
rect -90 982 -60 1182
rect 62 982 92 1182
rect 214 982 244 1784
rect 366 1584 396 1784
rect 366 982 396 1182
<< ndiff >>
rect -190 832 -90 862
rect -190 90 -160 832
rect -120 90 -90 832
rect -190 60 -90 90
rect -60 832 62 862
rect -60 692 -32 832
rect 8 692 62 832
rect -60 662 62 692
rect 92 832 214 862
rect 92 692 146 832
rect 186 692 214 832
rect 92 662 214 692
rect 244 830 366 862
rect 244 690 296 830
rect 336 690 366 830
rect 244 662 366 690
rect 396 832 492 862
rect 396 692 424 832
rect 464 692 492 832
rect 396 662 492 692
rect -60 260 -10 662
rect -60 230 62 260
rect -60 90 -32 230
rect 8 90 62 230
rect -60 60 62 90
rect 92 230 214 260
rect 92 90 146 230
rect 186 90 214 230
rect 92 60 214 90
rect 244 228 346 260
rect 244 88 276 228
rect 316 88 346 228
rect 244 60 346 88
rect 376 230 472 260
rect 376 90 404 230
rect 444 90 472 230
rect 376 60 472 90
<< pdiff >>
rect -190 1756 -90 1784
rect -190 1616 -160 1756
rect -120 1616 -90 1756
rect -190 1584 -90 1616
rect -60 1756 42 1784
rect -60 1616 -28 1756
rect 12 1616 42 1756
rect -60 1584 42 1616
rect 72 1754 214 1784
rect 72 1614 120 1754
rect 160 1614 214 1754
rect 72 1584 214 1614
rect 164 1182 214 1584
rect -190 1154 -90 1182
rect -190 1014 -160 1154
rect -120 1014 -90 1154
rect -190 982 -90 1014
rect -60 1154 62 1182
rect -60 1014 -8 1154
rect 32 1014 62 1154
rect -60 982 62 1014
rect 92 1152 214 1182
rect 92 1012 120 1152
rect 160 1012 214 1152
rect 92 982 214 1012
rect 244 1754 366 1784
rect 244 1614 272 1754
rect 312 1614 366 1754
rect 244 1584 366 1614
rect 396 1754 518 1784
rect 396 1614 450 1754
rect 490 1614 518 1754
rect 396 1584 518 1614
rect 244 1182 294 1584
rect 244 1152 366 1182
rect 244 1012 272 1152
rect 312 1012 366 1152
rect 244 982 366 1012
rect 396 1152 518 1182
rect 396 1012 450 1152
rect 490 1012 518 1152
rect 396 982 518 1012
<< ndiffc >>
rect -160 90 -120 832
rect -32 692 8 832
rect 146 692 186 832
rect 296 690 336 830
rect 424 692 464 832
rect -32 90 8 230
rect 146 90 186 230
rect 276 88 316 228
rect 404 90 444 230
<< pdiffc >>
rect -160 1616 -120 1756
rect -28 1616 12 1756
rect 120 1614 160 1754
rect -160 1014 -120 1154
rect -8 1014 32 1154
rect 120 1012 160 1152
rect 272 1614 312 1754
rect 450 1614 490 1754
rect 272 1012 312 1152
rect 450 1012 490 1152
<< psubdiff >>
rect 274 -22 474 6
rect 274 -62 304 -22
rect 444 -62 474 -22
rect 274 -90 474 -62
<< nsubdiff >>
rect -26 1910 174 1940
rect -26 1870 4 1910
rect 144 1870 174 1910
rect -26 1840 174 1870
<< psubdiffcont >>
rect 304 -62 444 -22
<< nsubdiffcont >>
rect 4 1870 144 1910
<< poly >>
rect -90 1784 -60 1812
rect 42 1784 72 1810
rect 214 1784 244 1810
rect 366 1784 396 1810
rect -90 1564 -60 1584
rect -156 1532 -60 1564
rect -156 1238 -126 1532
rect 42 1502 72 1584
rect 20 1476 110 1502
rect 20 1436 46 1476
rect 86 1436 110 1476
rect 20 1412 110 1436
rect -84 1344 6 1370
rect -84 1304 -58 1344
rect -18 1310 6 1344
rect -18 1304 12 1310
rect -84 1280 12 1304
rect -18 1238 12 1280
rect -156 1208 -60 1238
rect -18 1208 92 1238
rect -90 1182 -60 1208
rect 62 1182 92 1208
rect 366 1560 396 1584
rect 318 1536 408 1560
rect 318 1496 342 1536
rect 382 1496 408 1536
rect 318 1470 408 1496
rect 388 1404 478 1428
rect 388 1364 412 1404
rect 452 1364 478 1404
rect 388 1338 478 1364
rect 388 1308 418 1338
rect 366 1278 418 1308
rect 366 1182 396 1278
rect -90 862 -60 982
rect 62 862 92 982
rect 214 862 244 982
rect 366 862 396 982
rect 62 566 92 662
rect 62 536 104 566
rect 74 506 104 536
rect 74 480 164 506
rect 74 440 98 480
rect 138 440 164 480
rect 74 416 164 440
rect 6 348 96 374
rect 6 308 30 348
rect 70 308 96 348
rect 6 284 96 308
rect 62 260 92 284
rect 214 260 244 662
rect 366 642 396 662
rect 366 612 448 642
rect 286 546 376 570
rect 286 506 312 546
rect 352 506 376 546
rect 286 480 376 506
rect 286 306 316 480
rect 418 438 448 612
rect 359 414 449 438
rect 359 374 385 414
rect 425 374 449 414
rect 359 348 449 374
rect 286 276 376 306
rect 346 260 376 276
rect -90 24 -60 60
rect 62 34 92 60
rect 214 24 244 60
rect 346 34 376 60
rect -150 -2 -60 24
rect -150 -42 -126 -2
rect -86 -42 -60 -2
rect -150 -66 -60 -42
rect 154 -2 244 24
rect 154 -42 180 -2
rect 220 -42 244 -2
rect 154 -66 244 -42
<< polycont >>
rect 46 1436 86 1476
rect -58 1304 -18 1344
rect 342 1496 382 1536
rect 412 1364 452 1404
rect 98 440 138 480
rect 30 308 70 348
rect 312 506 352 546
rect 385 374 425 414
rect -126 -42 -86 -2
rect 180 -42 220 -2
<< locali >>
rect -16 1910 164 1930
rect -16 1870 4 1910
rect 144 1870 164 1910
rect -16 1850 164 1870
rect 100 1774 134 1850
rect -182 1756 -100 1774
rect -182 1628 -160 1756
rect -226 1616 -160 1628
rect -120 1616 -100 1756
rect -226 1594 -100 1616
rect -50 1756 32 1774
rect -50 1616 -28 1756
rect 12 1616 32 1756
rect -50 1594 32 1616
rect 100 1754 180 1774
rect 100 1614 120 1754
rect 160 1614 180 1754
rect 100 1594 180 1614
rect 252 1754 332 1774
rect 252 1614 272 1754
rect 312 1614 332 1754
rect 252 1594 332 1614
rect 430 1754 510 1774
rect 430 1614 450 1754
rect 490 1628 510 1754
rect 490 1614 556 1628
rect 430 1594 556 1614
rect -50 1554 -16 1594
rect -84 1520 -16 1554
rect -84 1370 -50 1520
rect 20 1476 110 1502
rect 20 1436 46 1476
rect 86 1436 110 1476
rect 20 1412 110 1436
rect -84 1344 6 1370
rect -84 1304 -58 1344
rect -18 1304 6 1344
rect -84 1280 6 1304
rect 76 1240 110 1412
rect 12 1206 110 1240
rect 12 1172 46 1206
rect 146 1172 180 1594
rect 318 1536 408 1560
rect 318 1504 342 1536
rect 310 1496 342 1504
rect 382 1496 408 1536
rect 310 1470 408 1496
rect 310 1266 344 1470
rect 442 1428 476 1594
rect 388 1404 478 1428
rect 388 1364 412 1404
rect 452 1364 478 1404
rect 388 1338 478 1364
rect 310 1232 464 1266
rect 430 1172 464 1232
rect -226 1154 -100 1172
rect -226 1138 -160 1154
rect -182 1014 -160 1138
rect -120 1014 -100 1154
rect -182 992 -100 1014
rect -30 1154 52 1172
rect -30 1014 -8 1154
rect 32 1014 52 1154
rect -30 992 52 1014
rect 100 1152 180 1172
rect 100 1012 120 1152
rect 160 1012 180 1152
rect 100 992 180 1012
rect 252 1152 332 1172
rect 252 1012 272 1152
rect 312 1012 332 1152
rect 18 956 52 992
rect 252 990 332 1012
rect 430 1152 556 1172
rect 430 1012 450 1152
rect 490 1138 556 1152
rect 490 1012 510 1138
rect 430 992 510 1012
rect 18 922 160 956
rect 430 922 464 992
rect -180 832 -100 854
rect -180 90 -160 832
rect -120 90 -100 832
rect -52 832 28 854
rect -52 692 -32 832
rect 8 692 28 832
rect -52 672 28 692
rect 126 852 160 922
rect 322 888 464 922
rect 322 852 356 888
rect 126 832 206 852
rect 126 692 146 832
rect 186 692 206 832
rect 126 672 206 692
rect 274 830 356 852
rect 274 690 296 830
rect 336 690 356 830
rect 274 672 356 690
rect 404 832 484 852
rect 404 692 424 832
rect 464 692 484 832
rect 404 672 484 692
rect 126 612 160 672
rect 6 578 160 612
rect 6 374 40 578
rect 286 570 320 672
rect 286 546 376 570
rect 286 506 312 546
rect 352 506 376 546
rect 74 480 164 506
rect 286 480 376 506
rect 450 506 484 672
rect 74 440 98 480
rect 138 440 164 480
rect 450 472 518 506
rect 74 416 164 440
rect 6 348 96 374
rect 6 308 30 348
rect 70 308 96 348
rect 6 284 96 308
rect 130 250 164 416
rect 359 414 449 438
rect 359 382 385 414
rect 302 374 385 382
rect 425 374 449 414
rect 302 348 449 374
rect 302 250 336 348
rect 484 314 518 472
rect 430 280 518 314
rect 430 250 464 280
rect -180 70 -100 90
rect -52 230 28 250
rect -52 90 -32 230
rect 8 90 28 230
rect -52 70 28 90
rect 126 230 206 250
rect 126 90 146 230
rect 186 90 206 230
rect 126 70 206 90
rect 254 228 336 250
rect 254 88 276 228
rect 316 88 336 228
rect 254 70 336 88
rect 384 230 464 250
rect 384 90 404 230
rect 444 90 464 230
rect 384 70 464 90
rect -150 -2 -60 24
rect -150 -42 -126 -2
rect -86 -42 -60 -2
rect -150 -66 -60 -42
rect 154 -2 244 24
rect 384 -2 418 70
rect 154 -42 180 -2
rect 220 -42 244 -2
rect 154 -66 244 -42
rect -150 -144 -116 -66
rect 210 -144 244 -66
rect 284 -22 464 -2
rect 284 -62 304 -22
rect 444 -62 464 -22
rect 284 -82 464 -62
rect -150 -152 -98 -144
rect -150 -186 -142 -152
rect -106 -186 -98 -152
rect -150 -194 -98 -186
rect 192 -152 244 -144
rect 192 -186 200 -152
rect 236 -186 244 -152
rect 192 -194 244 -186
<< viali >>
rect 4 1870 144 1910
rect 120 1614 160 1754
rect 120 1012 160 1152
rect -160 90 -120 832
rect 424 692 464 832
rect 404 90 444 230
rect 304 -62 444 -22
rect -142 -186 -106 -152
rect 200 -186 236 -152
<< metal1 >>
rect -226 1910 556 1930
rect -226 1870 4 1910
rect 144 1870 556 1910
rect -226 1754 556 1870
rect -226 1614 120 1754
rect 160 1614 556 1754
rect -226 1152 556 1614
rect -226 1012 120 1152
rect 160 1012 556 1152
rect -226 994 556 1012
rect -226 852 484 854
rect -226 832 556 852
rect -226 90 -160 832
rect -120 692 424 832
rect 464 692 556 832
rect -120 230 556 692
rect -120 90 404 230
rect 444 90 556 230
rect -226 -22 556 90
rect -226 -62 304 -22
rect 444 -62 556 -22
rect -226 -86 556 -62
rect -226 -152 556 -144
rect -226 -186 -142 -152
rect -106 -186 200 -152
rect 236 -186 556 -152
rect -226 -194 556 -186
<< labels >>
rlabel metal1 -226 1850 -226 1850 7 VP
port 1 w
rlabel metal1 -226 -170 -226 -170 7 CLK
port 5 w
rlabel metal1 -226 402 -226 402 7 VN
port 4 w
rlabel locali -226 1610 -226 1610 7 D
port 2 w
rlabel locali -226 1154 -226 1154 7 Dbar
port 3 w
rlabel locali 556 1612 556 1612 3 Q
port 6 e
rlabel locali 556 1156 556 1156 3 Qbar
port 7 e
<< end >>
