magic
tech sky130A
magscale 1 2
timestamp 1695950478
<< nwell >>
rect -414 1142 -4 1422
<< nmos >>
rect -174 863 -144 1063
<< pmos >>
rect -174 1182 -144 1382
<< ndiff >>
rect -274 1033 -174 1063
rect -274 893 -244 1033
rect -204 893 -174 1033
rect -274 863 -174 893
rect -144 1033 -44 1063
rect -144 893 -114 1033
rect -74 893 -44 1033
rect -144 863 -44 893
<< pdiff >>
rect -274 1352 -174 1382
rect -274 1212 -244 1352
rect -204 1212 -174 1352
rect -274 1182 -174 1212
rect -144 1352 -44 1382
rect -144 1212 -114 1352
rect -74 1212 -44 1352
rect -144 1182 -44 1212
<< ndiffc >>
rect -244 893 -204 1033
rect -114 893 -74 1033
<< pdiffc >>
rect -244 1212 -204 1352
rect -114 1212 -74 1352
<< psubdiff >>
rect -374 1033 -274 1063
rect -374 893 -344 1033
rect -304 893 -274 1033
rect -374 863 -274 893
<< nsubdiff >>
rect -374 1352 -274 1382
rect -374 1212 -344 1352
rect -304 1212 -274 1352
rect -374 1182 -274 1212
<< psubdiffcont >>
rect -344 893 -304 1033
<< nsubdiffcont >>
rect -344 1212 -304 1352
<< poly >>
rect -174 1472 -94 1492
rect -174 1432 -154 1472
rect -114 1432 -94 1472
rect -174 1412 -94 1432
rect -174 1382 -144 1412
rect -174 1063 -144 1182
rect -174 833 -144 863
<< polycont >>
rect -154 1432 -114 1472
<< locali >>
rect -128 1792 -4 1826
rect -128 1492 -94 1792
rect -174 1472 -94 1492
rect -174 1432 -154 1472
rect -114 1432 -94 1472
rect -174 1412 -94 1432
rect -364 1352 -184 1372
rect -364 1212 -344 1352
rect -304 1212 -244 1352
rect -204 1212 -184 1352
rect -364 1192 -184 1212
rect -134 1370 -54 1372
rect -134 1352 -2 1370
rect -134 1212 -114 1352
rect -74 1336 -2 1352
rect -74 1212 -54 1336
rect -134 1192 -54 1212
rect -94 1053 -54 1192
rect -364 1033 -184 1053
rect -364 893 -344 1033
rect -304 893 -244 1033
rect -204 893 -184 1033
rect -364 873 -184 893
rect -134 1033 -54 1053
rect -134 893 -114 1033
rect -74 893 -54 1033
rect -134 873 -54 893
<< viali >>
rect -344 1212 -304 1352
rect -244 1212 -204 1352
rect -344 893 -304 1033
rect -244 893 -204 1033
<< metal1 >>
rect -414 1352 -4 1372
rect -414 1212 -344 1352
rect -304 1212 -244 1352
rect -204 1212 -4 1352
rect -414 1192 -4 1212
rect -414 1033 -4 1053
rect -414 893 -344 1033
rect -304 893 -244 1033
rect -204 893 -4 1033
rect -414 873 -4 893
use latch  latch_0
timestamp 1695946031
transform 1 0 222 0 1 198
box -226 -194 556 1978
use latch  latch_1
timestamp 1695946031
transform 1 0 1004 0 1 198
box -226 -194 556 1978
use latch  latch_2
timestamp 1695946031
transform 1 0 1786 0 1 198
box -226 -194 556 1978
use latch  latch_3
timestamp 1695946031
transform 1 0 2568 0 1 198
box -226 -194 556 1978
<< labels >>
rlabel metal1 -414 1282 -414 1282 7 VP
port 3 w
rlabel metal1 -414 963 -414 963 7 VN
port 4 w
<< end >>
