magic
tech sky130A
timestamp 1697505651
<< nwell >>
rect -148 6873 338 8266
rect -140 2157 346 3550
<< nmos >>
rect -80 8384 -30 9584
rect 20 8384 70 9584
rect 120 8384 170 9584
rect 220 8384 270 9584
rect 20 5639 70 6839
rect 120 5639 170 6839
rect -97 5434 303 5484
rect -97 5334 303 5384
rect -97 5234 303 5284
rect -97 5134 303 5184
rect -97 5034 303 5084
rect -97 4934 303 4984
rect 28 3584 78 4784
rect 128 3584 178 4784
rect -72 839 -22 2039
rect 28 839 78 2039
rect 128 839 178 2039
rect 228 839 278 2039
<< pmos >>
rect -80 6971 -30 8171
rect 20 6971 70 8171
rect 120 6971 170 8171
rect 220 6971 270 8171
rect -72 2252 -22 3452
rect 28 2252 78 3452
rect 128 2252 178 3452
rect 228 2252 278 3452
<< ndiff >>
rect -130 9570 -80 9584
rect -130 8398 -117 9570
rect -93 8398 -80 9570
rect -130 8384 -80 8398
rect -30 9570 20 9584
rect -30 8398 -17 9570
rect 7 8398 20 9570
rect -30 8384 20 8398
rect 70 9570 120 9584
rect 70 8398 83 9570
rect 107 8398 120 9570
rect 70 8384 120 8398
rect 170 9570 220 9584
rect 170 8398 183 9570
rect 207 8398 220 9570
rect 170 8384 220 8398
rect 270 9570 320 9584
rect 270 8398 283 9570
rect 307 8398 320 9570
rect 270 8384 320 8398
rect -30 6825 20 6839
rect -30 5653 -17 6825
rect 7 5653 20 6825
rect -30 5639 20 5653
rect 70 6825 120 6839
rect 70 5653 83 6825
rect 107 5653 120 6825
rect 70 5639 120 5653
rect 170 6825 220 6839
rect 170 5653 183 6825
rect 207 5653 220 6825
rect 170 5639 220 5653
rect -97 5520 303 5534
rect -97 5499 -82 5520
rect 289 5499 303 5520
rect -97 5484 303 5499
rect -97 5420 303 5434
rect -97 5399 -82 5420
rect 289 5399 303 5420
rect -97 5384 303 5399
rect -97 5320 303 5334
rect -97 5299 -82 5320
rect 289 5299 303 5320
rect -97 5284 303 5299
rect -97 5220 303 5234
rect -97 5199 -82 5220
rect 289 5199 303 5220
rect -97 5184 303 5199
rect -97 5120 303 5134
rect -97 5099 -82 5120
rect 289 5099 303 5120
rect -97 5084 303 5099
rect -97 5020 303 5034
rect -97 4999 -82 5020
rect 289 4999 303 5020
rect -97 4984 303 4999
rect -97 4920 303 4934
rect -97 4899 -82 4920
rect 289 4899 303 4920
rect -97 4884 303 4899
rect -22 4770 28 4784
rect -22 3598 -9 4770
rect 15 3598 28 4770
rect -22 3584 28 3598
rect 78 4770 128 4784
rect 78 3598 91 4770
rect 115 3598 128 4770
rect 78 3584 128 3598
rect 178 4770 228 4784
rect 178 3598 191 4770
rect 215 3598 228 4770
rect 178 3584 228 3598
rect -122 2025 -72 2039
rect -122 853 -109 2025
rect -85 853 -72 2025
rect -122 839 -72 853
rect -22 2025 28 2039
rect -22 853 -9 2025
rect 15 853 28 2025
rect -22 839 28 853
rect 78 2025 128 2039
rect 78 853 91 2025
rect 115 853 128 2025
rect 78 839 128 853
rect 178 2025 228 2039
rect 178 853 191 2025
rect 215 853 228 2025
rect 178 839 228 853
rect 278 2025 328 2039
rect 278 853 291 2025
rect 315 853 328 2025
rect 278 839 328 853
<< pdiff >>
rect -130 8157 -80 8171
rect -130 6985 -117 8157
rect -93 6985 -80 8157
rect -130 6971 -80 6985
rect -30 8157 20 8171
rect -30 6985 -17 8157
rect 7 6985 20 8157
rect -30 6971 20 6985
rect 70 8157 120 8171
rect 70 6985 83 8157
rect 107 6985 120 8157
rect 70 6971 120 6985
rect 170 8157 220 8171
rect 170 6985 183 8157
rect 207 6985 220 8157
rect 170 6971 220 6985
rect 270 8157 320 8171
rect 270 6985 283 8157
rect 307 6985 320 8157
rect 270 6971 320 6985
rect -122 3438 -72 3452
rect -122 2266 -109 3438
rect -85 2266 -72 3438
rect -122 2252 -72 2266
rect -22 3438 28 3452
rect -22 2266 -9 3438
rect 15 2266 28 3438
rect -22 2252 28 2266
rect 78 3438 128 3452
rect 78 2266 91 3438
rect 115 2266 128 3438
rect 78 2252 128 2266
rect 178 3438 228 3452
rect 178 2266 191 3438
rect 215 2266 228 3438
rect 178 2252 228 2266
rect 278 3438 328 3452
rect 278 2266 291 3438
rect 315 2266 328 3438
rect 278 2252 328 2266
<< ndiffc >>
rect -117 8398 -93 9570
rect -17 8398 7 9570
rect 83 8398 107 9570
rect 183 8398 207 9570
rect 283 8398 307 9570
rect -17 5653 7 6825
rect 83 5653 107 6825
rect 183 5653 207 6825
rect -82 5499 289 5520
rect -82 5399 289 5420
rect -82 5299 289 5320
rect -82 5199 289 5220
rect -82 5099 289 5120
rect -82 4999 289 5020
rect -82 4899 289 4920
rect -9 3598 15 4770
rect 91 3598 115 4770
rect 191 3598 215 4770
rect -109 853 -85 2025
rect -9 853 15 2025
rect 91 853 115 2025
rect 191 853 215 2025
rect 291 853 315 2025
<< pdiffc >>
rect -117 6985 -93 8157
rect -17 6985 7 8157
rect 83 6985 107 8157
rect 183 6985 207 8157
rect 283 6985 307 8157
rect -109 2266 -85 3438
rect -9 2266 15 3438
rect 91 2266 115 3438
rect 191 2266 215 3438
rect 291 2266 315 3438
<< psubdiff >>
rect 46 9647 148 9661
rect 46 9625 62 9647
rect 133 9625 148 9647
rect 46 9611 148 9625
rect 46 8315 148 8329
rect 46 8293 62 8315
rect 133 8293 148 8315
rect 46 8279 148 8293
rect -191 5243 -141 5257
rect -191 5172 -177 5243
rect -155 5172 -141 5243
rect -191 5157 -141 5172
rect 341 5242 391 5257
rect 341 5171 356 5242
rect 378 5171 391 5242
rect 341 5157 391 5171
rect 50 2130 152 2144
rect 50 2108 65 2130
rect 136 2108 152 2130
rect 50 2094 152 2108
rect 50 798 152 812
rect 50 776 65 798
rect 136 776 152 798
rect 50 762 152 776
<< nsubdiff >>
rect 46 8234 148 8248
rect 46 8212 62 8234
rect 133 8212 148 8234
rect 46 8198 148 8212
rect 46 6928 148 6942
rect 46 6906 62 6928
rect 133 6906 148 6928
rect 46 6892 148 6906
rect 50 3517 152 3531
rect 50 3495 65 3517
rect 136 3495 152 3517
rect 50 3481 152 3495
rect 50 2211 152 2225
rect 50 2189 65 2211
rect 136 2189 152 2211
rect 50 2175 152 2189
<< psubdiffcont >>
rect 62 9625 133 9647
rect 62 8293 133 8315
rect -177 5172 -155 5243
rect 356 5171 378 5242
rect 65 2108 136 2130
rect 65 776 136 798
<< nsubdiffcont >>
rect 62 8212 133 8234
rect 62 6906 133 6928
rect 65 3495 136 3517
rect 65 2189 136 2211
<< poly >>
rect -224 9669 270 9684
rect -80 9584 -30 9669
rect 20 9584 70 9597
rect 120 9584 170 9597
rect 220 9584 270 9669
rect -80 8371 -30 8384
rect 20 8376 70 8384
rect 120 8376 170 8384
rect 20 8350 170 8376
rect 220 8371 270 8384
rect 20 8342 314 8350
rect 20 8335 285 8342
rect 276 8320 285 8335
rect 306 8320 314 8342
rect 276 8312 314 8320
rect -224 8256 270 8271
rect -80 8171 -30 8256
rect 20 8171 70 8184
rect 120 8171 170 8184
rect 220 8171 270 8256
rect -80 6958 -30 6971
rect 20 6963 70 6971
rect 120 6963 170 6971
rect 20 6948 170 6963
rect 220 6958 270 6971
rect 20 6933 40 6948
rect -224 6918 40 6933
rect 20 6839 70 6852
rect 120 6839 170 6852
rect -81 5641 -43 5649
rect -81 5619 -73 5641
rect -52 5626 -43 5641
rect 20 5626 70 5639
rect -52 5619 70 5626
rect -81 5611 70 5619
rect 120 5590 170 5639
rect -75 5582 170 5590
rect -75 5560 -67 5582
rect -46 5575 170 5582
rect -46 5560 -37 5575
rect -75 5552 -37 5560
rect -127 5434 -97 5484
rect 303 5434 333 5484
rect -127 5384 -112 5434
rect 318 5384 333 5434
rect -224 5364 -186 5372
rect -224 5342 -216 5364
rect -195 5342 -186 5364
rect -224 5334 -186 5342
rect -127 5334 -97 5384
rect 303 5334 333 5384
rect -224 5139 -209 5334
rect -186 5305 -148 5313
rect -186 5283 -178 5305
rect -157 5283 -148 5305
rect -186 5275 -148 5283
rect -127 5284 -112 5334
rect 318 5284 333 5334
rect -127 5234 -97 5284
rect 303 5234 333 5284
rect -127 5184 -112 5234
rect 318 5184 333 5234
rect -224 5131 -148 5139
rect -224 5124 -178 5131
rect -186 5109 -178 5124
rect -157 5109 -148 5131
rect -186 5101 -148 5109
rect -127 5134 -97 5184
rect 303 5134 333 5184
rect -127 5084 -112 5134
rect 318 5084 333 5134
rect -127 5034 -97 5084
rect 303 5034 333 5084
rect -127 4984 -112 5034
rect 318 4984 333 5034
rect -127 4949 -97 4984
rect -224 4934 -97 4949
rect 303 4934 333 4984
rect -67 4858 -29 4866
rect -67 4836 -59 4858
rect -38 4843 -29 4858
rect -38 4836 178 4843
rect -67 4828 178 4836
rect -74 4799 78 4807
rect -74 4777 -66 4799
rect -45 4792 78 4799
rect -45 4777 -36 4792
rect 28 4784 78 4792
rect 128 4784 178 4828
rect -74 4769 -36 4777
rect 28 3571 78 3584
rect 128 3571 178 3584
rect -224 3486 44 3501
rect 28 3475 44 3486
rect -72 3452 -22 3465
rect 28 3460 178 3475
rect 28 3452 78 3460
rect 128 3452 178 3460
rect 228 3452 278 3465
rect -72 2167 -22 2252
rect 28 2239 78 2252
rect 128 2239 178 2252
rect 228 2167 278 2252
rect -224 2152 278 2167
rect -116 2103 -78 2111
rect -116 2081 -108 2103
rect -87 2088 -78 2103
rect -87 2081 178 2088
rect -116 2073 178 2081
rect -72 2039 -22 2052
rect 28 2047 178 2073
rect 28 2039 78 2047
rect 128 2039 178 2047
rect 228 2039 278 2052
rect -72 754 -22 839
rect 28 826 78 839
rect 128 826 178 839
rect 228 754 278 839
rect -224 739 278 754
<< polycont >>
rect 285 8320 306 8342
rect -73 5619 -52 5641
rect -67 5560 -46 5582
rect -216 5342 -195 5364
rect -178 5283 -157 5305
rect -178 5109 -157 5131
rect -59 4836 -38 4858
rect -66 4777 -45 4799
rect -108 2081 -87 2103
<< locali >>
rect 52 9647 142 9656
rect 52 9625 62 9647
rect 133 9625 142 9647
rect 52 9616 142 9625
rect -124 9570 -86 9578
rect -124 8398 -117 9570
rect -93 8398 -86 9570
rect -124 8157 -86 8398
rect -24 9570 14 9578
rect -24 8398 -17 9570
rect 7 8398 14 9570
rect -24 8390 14 8398
rect 76 9570 114 9616
rect 76 8398 83 9570
rect 107 8398 114 9570
rect 76 8324 114 8398
rect 176 9570 214 9578
rect 176 8398 183 9570
rect 207 8398 214 9570
rect 176 8390 214 8398
rect 276 9570 314 9578
rect 276 8398 283 9570
rect 307 8398 314 9570
rect 276 8342 314 8398
rect 52 8315 142 8324
rect 52 8293 62 8315
rect 133 8293 142 8315
rect 52 8284 142 8293
rect 276 8320 285 8342
rect 306 8320 314 8342
rect 52 8234 142 8243
rect 52 8212 62 8234
rect 133 8212 142 8234
rect 52 8203 142 8212
rect -124 6985 -117 8157
rect -93 6985 -86 8157
rect -124 6977 -86 6985
rect -24 8157 14 8165
rect -24 6985 -17 8157
rect 7 6985 14 8157
rect -24 6825 14 6985
rect 76 8157 114 8203
rect 76 6985 83 8157
rect 107 6985 114 8157
rect 76 6937 114 6985
rect 176 8157 214 8165
rect 176 6985 183 8157
rect 207 6985 214 8157
rect 52 6928 142 6937
rect 52 6906 62 6928
rect 133 6906 142 6928
rect 52 6897 142 6906
rect -24 5653 -17 6825
rect 7 5653 14 6825
rect -81 5641 -43 5649
rect -24 5645 14 5653
rect 76 6825 114 6839
rect 76 5653 83 6825
rect 107 5653 114 6825
rect -81 5628 -73 5641
rect -224 5619 -73 5628
rect -52 5619 -43 5641
rect -224 5611 -43 5619
rect -224 5372 -206 5611
rect -75 5582 -37 5590
rect -75 5569 -67 5582
rect -166 5560 -67 5569
rect -46 5560 -37 5582
rect -166 5552 -37 5560
rect -224 5364 -186 5372
rect -224 5342 -216 5364
rect -195 5342 -186 5364
rect -224 5334 -186 5342
rect -166 5313 -148 5552
rect 76 5528 114 5653
rect 176 6825 214 6985
rect 276 8157 314 8320
rect 276 6985 283 8157
rect 307 6985 314 8157
rect 276 6977 314 6985
rect 176 5653 183 6825
rect 207 5653 214 6825
rect 176 5645 214 5653
rect -186 5305 -148 5313
rect -186 5292 -178 5305
rect -224 5283 -178 5292
rect -157 5283 -148 5305
rect -124 5520 297 5528
rect -124 5499 -82 5520
rect 289 5499 297 5520
rect -124 5490 297 5499
rect -124 5328 -107 5490
rect -90 5420 331 5428
rect -90 5399 -82 5420
rect 289 5399 331 5420
rect -90 5390 331 5399
rect -124 5320 297 5328
rect -124 5299 -82 5320
rect 289 5299 297 5320
rect -124 5290 297 5299
rect -224 5275 -148 5283
rect -224 4807 -206 5275
rect -185 5243 -147 5251
rect -185 5172 -177 5243
rect -155 5228 -147 5243
rect 314 5228 331 5390
rect 348 5242 386 5250
rect 348 5228 356 5242
rect -155 5220 356 5228
rect -155 5199 -82 5220
rect 289 5199 356 5220
rect -155 5190 356 5199
rect -155 5172 -147 5190
rect -185 5163 -147 5172
rect -186 5131 -148 5139
rect -186 5109 -178 5131
rect -157 5109 -148 5131
rect -186 5101 -148 5109
rect -169 4866 -151 5101
rect -124 5028 -107 5190
rect 348 5171 356 5190
rect 378 5171 386 5242
rect 348 5163 386 5171
rect -90 5120 331 5128
rect -90 5099 -82 5120
rect 289 5099 331 5120
rect -90 5090 331 5099
rect -124 5020 297 5028
rect -124 4999 -82 5020
rect 289 4999 297 5020
rect -124 4990 297 4999
rect 314 4928 331 5090
rect -90 4920 331 4928
rect -90 4899 -82 4920
rect 289 4899 331 4920
rect -90 4890 331 4899
rect -169 4858 -29 4866
rect -169 4849 -59 4858
rect -67 4836 -59 4849
rect -38 4836 -29 4858
rect -67 4828 -29 4836
rect -224 4799 -36 4807
rect -224 4790 -66 4799
rect -74 4777 -66 4790
rect -45 4777 -36 4799
rect -74 4769 -36 4777
rect -16 4770 22 4778
rect -16 3598 -9 4770
rect 15 3598 22 4770
rect -116 3438 -78 3446
rect -116 2266 -109 3438
rect -85 2266 -78 3438
rect -116 2103 -78 2266
rect -16 3438 22 3598
rect 84 4770 122 4890
rect 84 3598 91 4770
rect 115 3598 122 4770
rect 84 3584 122 3598
rect 184 4770 222 4778
rect 184 3598 191 4770
rect 215 3598 222 4770
rect 56 3517 146 3526
rect 56 3495 65 3517
rect 136 3495 146 3517
rect 56 3486 146 3495
rect -16 2266 -9 3438
rect 15 2266 22 3438
rect -16 2258 22 2266
rect 84 3438 122 3486
rect 84 2266 91 3438
rect 115 2266 122 3438
rect 84 2220 122 2266
rect 184 3438 222 3598
rect 184 2266 191 3438
rect 215 2266 222 3438
rect 184 2258 222 2266
rect 284 3438 457 3446
rect 284 2266 291 3438
rect 315 3429 457 3438
rect 315 2266 322 3429
rect 56 2211 146 2220
rect 56 2189 65 2211
rect 136 2189 146 2211
rect 56 2180 146 2189
rect -116 2081 -108 2103
rect -87 2081 -78 2103
rect 56 2130 146 2139
rect 56 2108 65 2130
rect 136 2108 146 2130
rect 56 2099 146 2108
rect -116 2025 -78 2081
rect -116 853 -109 2025
rect -85 853 -78 2025
rect -116 845 -78 853
rect -16 2025 22 2033
rect -16 853 -9 2025
rect 15 853 22 2025
rect -16 845 22 853
rect 84 2025 122 2099
rect 84 853 91 2025
rect 115 853 122 2025
rect 84 807 122 853
rect 184 2025 222 2033
rect 184 853 191 2025
rect 215 853 222 2025
rect 184 845 222 853
rect 284 2025 322 2266
rect 284 853 291 2025
rect 315 853 322 2025
rect 284 845 322 853
rect 56 798 146 807
rect 56 776 65 798
rect 136 776 146 798
rect 56 767 146 776
<< viali >>
rect 62 9625 133 9647
rect 62 8293 133 8315
rect 62 8212 133 8234
rect 62 6906 133 6928
rect -177 5172 -155 5243
rect 356 5171 378 5242
rect 65 3495 136 3517
rect 65 2189 136 2211
rect 65 2108 136 2130
rect 65 776 136 798
<< metal1 >>
rect -122 9647 148 9670
rect -122 9625 62 9647
rect 133 9625 148 9647
rect -122 9610 148 9625
rect -122 8380 20 9610
rect -122 8315 148 8380
rect -122 8293 62 8315
rect 133 8293 148 8315
rect -122 8278 148 8293
rect -122 7341 20 8278
rect 201 8248 344 9684
rect 46 8234 344 8248
rect 46 8212 62 8234
rect 133 8212 344 8234
rect 46 8198 344 8212
rect -123 5257 19 7341
rect 201 6942 344 8198
rect 46 6928 344 6942
rect 46 6906 62 6928
rect 133 6906 344 6928
rect 46 6892 344 6906
rect 201 5334 344 6892
rect 201 5275 457 5334
rect -191 5243 391 5257
rect -191 5172 -177 5243
rect -155 5242 391 5243
rect -155 5172 356 5242
rect -191 5171 356 5172
rect 378 5171 391 5242
rect -191 5157 391 5171
rect -123 4715 19 5157
rect 412 5132 457 5275
rect -122 2140 19 4715
rect 201 5072 457 5132
rect 201 4803 344 5072
rect 201 3531 342 4803
rect 50 3517 342 3531
rect 50 3495 65 3517
rect 136 3495 342 3517
rect 50 3481 342 3495
rect 201 2709 342 3481
rect 201 2225 343 2709
rect 50 2211 343 2225
rect 50 2189 65 2211
rect 136 2189 343 2211
rect 50 2175 343 2189
rect -122 2130 153 2140
rect -122 2108 65 2130
rect 136 2108 153 2130
rect -122 2094 153 2108
rect -122 813 50 2094
rect 201 1455 343 2175
rect -122 798 153 813
rect -122 776 65 798
rect 136 776 153 798
rect -122 739 153 776
rect 201 758 342 1455
<< labels >>
rlabel metal1 15 739 15 739 5 VN
port 11 s
rlabel metal1 276 9684 276 9684 1 VP
port 10 n
rlabel locali 457 3437 457 3437 3 Vout
port 12 e
rlabel poly -224 9676 -224 9676 7 VcnT
port 1 w
rlabel poly -224 8264 -224 8264 7 VcpT
port 2 w
rlabel poly -224 6925 -224 6925 7 VbpT
port 3 w
rlabel poly -224 4941 -224 4941 7 Vbn
port 6 w
rlabel locali -224 5284 -224 5284 7 V1
port 4 w
rlabel poly -224 5132 -224 5132 7 V2
port 5 w
rlabel poly -224 3493 -224 3493 7 Vbp
port 7 w
rlabel poly -224 2159 -224 2159 7 Vcp
port 8 w
rlabel poly -224 746 -224 746 7 Vcn
port 9 w
<< end >>
