magic
tech sky130A
timestamp 1697568761
<< nwell >>
rect -70 3990 1695 5320
rect 415 3900 535 3990
rect 1090 3900 1210 3990
rect 500 2570 620 2630
rect -70 1430 620 2570
rect 1005 2570 1125 2630
rect 1005 1430 1695 2570
rect -70 1310 700 1430
rect 925 1310 1695 1430
<< nmos >>
rect 0 2665 50 3865
rect 100 2665 150 3865
rect 200 2665 250 3865
rect 300 2665 350 3865
rect 400 2665 450 3865
rect 500 2665 550 3865
rect 735 2040 785 3240
rect 835 2040 885 3240
rect 1075 2665 1125 3865
rect 1175 2665 1225 3865
rect 1275 2665 1325 3865
rect 1375 2665 1425 3865
rect 1475 2665 1525 3865
rect 1575 2665 1625 3865
rect 0 0 50 1200
rect 100 0 150 1200
rect 200 0 250 1200
rect 300 0 350 1200
rect 400 0 450 1200
rect 500 0 550 1200
rect 735 0 785 1200
rect 835 0 885 1200
rect 1075 0 1125 1200
rect 1175 0 1225 1200
rect 1275 0 1325 1200
rect 1375 0 1425 1200
rect 1475 0 1525 1200
rect 1575 0 1625 1200
<< pmos >>
rect 0 4020 50 5220
rect 100 4020 150 5220
rect 200 4020 250 5220
rect 300 4020 350 5220
rect 400 4020 450 5220
rect 500 4020 550 5220
rect 735 4020 785 5220
rect 835 4020 885 5220
rect 1075 4020 1125 5220
rect 1175 4020 1225 5220
rect 1275 4020 1325 5220
rect 1375 4020 1425 5220
rect 1475 4020 1525 5220
rect 1575 4020 1625 5220
rect 0 1330 50 2530
rect 100 1330 150 2530
rect 200 1330 250 2530
rect 300 1330 350 2530
rect 400 1330 450 2530
rect 500 1330 550 2530
rect 1075 1330 1125 2530
rect 1175 1330 1225 2530
rect 1275 1330 1325 2530
rect 1375 1330 1425 2530
rect 1475 1330 1525 2530
rect 1575 1330 1625 2530
<< ndiff >>
rect -50 3845 0 3865
rect -50 2680 -35 3845
rect -15 2680 0 3845
rect -50 2665 0 2680
rect 50 3845 100 3865
rect 50 2680 65 3845
rect 85 2680 100 3845
rect 50 2665 100 2680
rect 150 3845 200 3865
rect 150 2680 165 3845
rect 185 2680 200 3845
rect 150 2665 200 2680
rect 250 3845 300 3865
rect 250 2680 265 3845
rect 285 2680 300 3845
rect 250 2665 300 2680
rect 350 3845 400 3865
rect 350 2680 365 3845
rect 385 2680 400 3845
rect 350 2665 400 2680
rect 450 3845 500 3865
rect 450 2680 465 3845
rect 485 2680 500 3845
rect 450 2665 500 2680
rect 550 3845 600 3865
rect 550 2680 565 3845
rect 585 2680 600 3845
rect 1025 3845 1075 3865
rect 550 2665 600 2680
rect 685 3220 735 3240
rect 685 2055 700 3220
rect 720 2055 735 3220
rect 685 2040 735 2055
rect 785 3220 835 3240
rect 785 2055 800 3220
rect 820 2055 835 3220
rect 785 2040 835 2055
rect 885 3220 935 3240
rect 885 2055 900 3220
rect 920 2055 935 3220
rect 1025 2680 1040 3845
rect 1060 2680 1075 3845
rect 1025 2665 1075 2680
rect 1125 3845 1175 3865
rect 1125 2680 1140 3845
rect 1160 2680 1175 3845
rect 1125 2665 1175 2680
rect 1225 3845 1275 3865
rect 1225 2680 1240 3845
rect 1260 2680 1275 3845
rect 1225 2665 1275 2680
rect 1325 3845 1375 3865
rect 1325 2680 1340 3845
rect 1360 2680 1375 3845
rect 1325 2665 1375 2680
rect 1425 3845 1475 3865
rect 1425 2680 1440 3845
rect 1460 2680 1475 3845
rect 1425 2665 1475 2680
rect 1525 3845 1575 3865
rect 1525 2680 1540 3845
rect 1560 2680 1575 3845
rect 1525 2665 1575 2680
rect 1625 3845 1675 3865
rect 1625 2680 1640 3845
rect 1660 2680 1675 3845
rect 1625 2665 1675 2680
rect 885 2040 935 2055
rect -50 1185 0 1200
rect -50 20 -35 1185
rect -15 20 0 1185
rect -50 0 0 20
rect 50 1185 100 1200
rect 50 20 65 1185
rect 85 20 100 1185
rect 50 0 100 20
rect 150 1185 200 1200
rect 150 20 165 1185
rect 185 20 200 1185
rect 150 0 200 20
rect 250 1185 300 1200
rect 250 20 265 1185
rect 285 20 300 1185
rect 250 0 300 20
rect 350 1185 400 1200
rect 350 20 365 1185
rect 385 20 400 1185
rect 350 0 400 20
rect 450 1185 500 1200
rect 450 20 465 1185
rect 485 20 500 1185
rect 450 0 500 20
rect 550 1185 600 1200
rect 550 20 565 1185
rect 585 20 600 1185
rect 550 0 600 20
rect 685 1180 735 1200
rect 685 15 700 1180
rect 720 15 735 1180
rect 685 0 735 15
rect 785 1180 835 1200
rect 785 15 800 1180
rect 820 15 835 1180
rect 785 0 835 15
rect 885 1180 935 1200
rect 885 15 900 1180
rect 920 15 935 1180
rect 885 0 935 15
rect 1025 1185 1075 1200
rect 1025 20 1040 1185
rect 1060 20 1075 1185
rect 1025 0 1075 20
rect 1125 1185 1175 1200
rect 1125 20 1140 1185
rect 1160 20 1175 1185
rect 1125 0 1175 20
rect 1225 1185 1275 1200
rect 1225 20 1240 1185
rect 1260 20 1275 1185
rect 1225 0 1275 20
rect 1325 1185 1375 1200
rect 1325 20 1340 1185
rect 1360 20 1375 1185
rect 1325 0 1375 20
rect 1425 1185 1475 1200
rect 1425 20 1440 1185
rect 1460 20 1475 1185
rect 1425 0 1475 20
rect 1525 1185 1575 1200
rect 1525 20 1540 1185
rect 1560 20 1575 1185
rect 1525 0 1575 20
rect 1625 1185 1675 1200
rect 1625 20 1640 1185
rect 1660 20 1675 1185
rect 1625 0 1675 20
<< pdiff >>
rect -50 5200 0 5220
rect -50 4035 -35 5200
rect -15 4035 0 5200
rect -50 4020 0 4035
rect 50 5200 100 5220
rect 50 4035 65 5200
rect 85 4035 100 5200
rect 50 4020 100 4035
rect 150 5200 200 5220
rect 150 4035 165 5200
rect 185 4035 200 5200
rect 150 4020 200 4035
rect 250 5200 300 5220
rect 250 4035 265 5200
rect 285 4035 300 5200
rect 250 4020 300 4035
rect 350 5200 400 5220
rect 350 4035 365 5200
rect 385 4035 400 5200
rect 350 4020 400 4035
rect 450 5200 500 5220
rect 450 4035 465 5200
rect 485 4035 500 5200
rect 450 4020 500 4035
rect 550 5200 600 5220
rect 550 4035 565 5200
rect 585 4035 600 5200
rect 550 4020 600 4035
rect 685 5200 735 5220
rect 685 4035 700 5200
rect 720 4035 735 5200
rect 685 4020 735 4035
rect 785 5200 835 5220
rect 785 4035 800 5200
rect 820 4035 835 5200
rect 785 4020 835 4035
rect 885 5200 935 5220
rect 885 4035 900 5200
rect 920 4035 935 5200
rect 885 4020 935 4035
rect 1025 5200 1075 5220
rect 1025 4035 1040 5200
rect 1060 4035 1075 5200
rect 1025 4020 1075 4035
rect 1125 5200 1175 5220
rect 1125 4035 1140 5200
rect 1160 4035 1175 5200
rect 1125 4020 1175 4035
rect 1225 5200 1275 5220
rect 1225 4035 1240 5200
rect 1260 4035 1275 5200
rect 1225 4020 1275 4035
rect 1325 5200 1375 5220
rect 1325 4035 1340 5200
rect 1360 4035 1375 5200
rect 1325 4020 1375 4035
rect 1425 5200 1475 5220
rect 1425 4035 1440 5200
rect 1460 4035 1475 5200
rect 1425 4020 1475 4035
rect 1525 5200 1575 5220
rect 1525 4035 1540 5200
rect 1560 4035 1575 5200
rect 1525 4020 1575 4035
rect 1625 5200 1675 5220
rect 1625 4035 1640 5200
rect 1660 4035 1675 5200
rect 1625 4020 1675 4035
rect -50 2515 0 2530
rect -50 1350 -35 2515
rect -15 1350 0 2515
rect -50 1330 0 1350
rect 50 2515 100 2530
rect 50 1350 65 2515
rect 85 1350 100 2515
rect 50 1330 100 1350
rect 150 2515 200 2530
rect 150 1350 165 2515
rect 185 1350 200 2515
rect 150 1330 200 1350
rect 250 2515 300 2530
rect 250 1350 265 2515
rect 285 1350 300 2515
rect 250 1330 300 1350
rect 350 2515 400 2530
rect 350 1350 365 2515
rect 385 1350 400 2515
rect 350 1330 400 1350
rect 450 2515 500 2530
rect 450 1350 465 2515
rect 485 1350 500 2515
rect 450 1330 500 1350
rect 550 2515 600 2530
rect 550 1350 565 2515
rect 585 1350 600 2515
rect 1025 2515 1075 2530
rect 550 1330 600 1350
rect 1025 1350 1040 2515
rect 1060 1350 1075 2515
rect 1025 1330 1075 1350
rect 1125 2515 1175 2530
rect 1125 1350 1140 2515
rect 1160 1350 1175 2515
rect 1125 1330 1175 1350
rect 1225 2515 1275 2530
rect 1225 1350 1240 2515
rect 1260 1350 1275 2515
rect 1225 1330 1275 1350
rect 1325 2515 1375 2530
rect 1325 1350 1340 2515
rect 1360 1350 1375 2515
rect 1325 1330 1375 1350
rect 1425 2515 1475 2530
rect 1425 1350 1440 2515
rect 1460 1350 1475 2515
rect 1425 1330 1475 1350
rect 1525 2515 1575 2530
rect 1525 1350 1540 2515
rect 1560 1350 1575 2515
rect 1525 1330 1575 1350
rect 1625 2515 1675 2530
rect 1625 1350 1640 2515
rect 1660 1350 1675 2515
rect 1625 1330 1675 1350
<< ndiffc >>
rect -35 2680 -15 3845
rect 65 2680 85 3845
rect 165 2680 185 3845
rect 265 2680 285 3845
rect 365 2680 385 3845
rect 465 2680 485 3845
rect 565 2680 585 3845
rect 700 2055 720 3220
rect 800 2055 820 3220
rect 900 2055 920 3220
rect 1040 2680 1060 3845
rect 1140 2680 1160 3845
rect 1240 2680 1260 3845
rect 1340 2680 1360 3845
rect 1440 2680 1460 3845
rect 1540 2680 1560 3845
rect 1640 2680 1660 3845
rect -35 20 -15 1185
rect 65 20 85 1185
rect 165 20 185 1185
rect 265 20 285 1185
rect 365 20 385 1185
rect 465 20 485 1185
rect 565 20 585 1185
rect 700 15 720 1180
rect 800 15 820 1180
rect 900 15 920 1180
rect 1040 20 1060 1185
rect 1140 20 1160 1185
rect 1240 20 1260 1185
rect 1340 20 1360 1185
rect 1440 20 1460 1185
rect 1540 20 1560 1185
rect 1640 20 1660 1185
<< pdiffc >>
rect -35 4035 -15 5200
rect 65 4035 85 5200
rect 165 4035 185 5200
rect 265 4035 285 5200
rect 365 4035 385 5200
rect 465 4035 485 5200
rect 565 4035 585 5200
rect 700 4035 720 5200
rect 800 4035 820 5200
rect 900 4035 920 5200
rect 1040 4035 1060 5200
rect 1140 4035 1160 5200
rect 1240 4035 1260 5200
rect 1340 4035 1360 5200
rect 1440 4035 1460 5200
rect 1540 4035 1560 5200
rect 1640 4035 1660 5200
rect -35 1350 -15 2515
rect 65 1350 85 2515
rect 165 1350 185 2515
rect 265 1350 285 2515
rect 365 1350 385 2515
rect 465 1350 485 2515
rect 565 1350 585 2515
rect 1040 1350 1060 2515
rect 1140 1350 1160 2515
rect 1240 1350 1260 2515
rect 1340 1350 1360 2515
rect 1440 1350 1460 2515
rect 1540 1350 1560 2515
rect 1640 1350 1660 2515
<< psubdiff >>
rect -130 3850 -80 3865
rect -130 3800 -115 3850
rect -95 3800 -80 3850
rect -130 3785 -80 3800
rect 635 3220 685 3240
rect -50 2620 30 2635
rect -50 2600 -35 2620
rect 15 2600 30 2620
rect -50 2585 30 2600
rect 635 2055 650 3220
rect 670 2055 685 3220
rect 635 2040 685 2055
rect 935 3220 985 3240
rect 935 2055 950 3220
rect 970 2055 985 3220
rect 1705 3850 1755 3865
rect 1705 3800 1720 3850
rect 1740 3800 1755 3850
rect 1705 3785 1755 3800
rect 1595 2620 1675 2635
rect 1595 2600 1610 2620
rect 1660 2600 1675 2620
rect 1595 2585 1675 2600
rect 935 2040 985 2055
rect 35 1275 115 1290
rect 35 1255 50 1275
rect 100 1255 115 1275
rect 35 1240 115 1255
rect 1510 1275 1590 1290
rect 1510 1255 1525 1275
rect 1575 1255 1590 1275
rect 1510 1240 1590 1255
rect 635 1180 685 1200
rect 635 15 650 1180
rect 670 15 685 1180
rect 635 0 685 15
rect 935 1180 985 1200
rect 935 15 950 1180
rect 970 15 985 1180
rect 935 0 985 15
rect 35 -45 115 -30
rect 35 -65 50 -45
rect 100 -65 115 -45
rect 35 -80 115 -65
rect 1510 -45 1590 -30
rect 1510 -65 1525 -45
rect 1575 -65 1590 -45
rect 1510 -80 1590 -65
<< nsubdiff >>
rect 435 5285 515 5300
rect 435 5265 450 5285
rect 500 5265 515 5285
rect 435 5250 515 5265
rect 1110 5285 1190 5300
rect 1110 5265 1125 5285
rect 1175 5265 1190 5285
rect 1110 5250 1190 5265
rect 635 5200 685 5220
rect 635 4035 650 5200
rect 670 4035 685 5200
rect 635 4020 685 4035
rect 935 5200 985 5220
rect 935 4035 950 5200
rect 970 4035 985 5200
rect 935 4020 985 4035
rect 435 3955 515 3970
rect 435 3935 450 3955
rect 500 3935 515 3955
rect 435 3920 515 3935
rect 1110 3955 1190 3970
rect 1110 3935 1125 3955
rect 1175 3935 1190 3955
rect 1110 3920 1190 3935
rect 520 2595 600 2610
rect 520 2575 535 2595
rect 585 2575 600 2595
rect 520 2560 600 2575
rect 1025 2595 1105 2610
rect 1025 2575 1040 2595
rect 1090 2575 1105 2595
rect 1025 2560 1105 2575
rect 630 1395 680 1410
rect 630 1345 645 1395
rect 665 1345 680 1395
rect 630 1330 680 1345
rect 945 1395 995 1410
rect 945 1345 960 1395
rect 980 1345 995 1395
rect 945 1330 995 1345
<< psubdiffcont >>
rect -115 3800 -95 3850
rect -35 2600 15 2620
rect 650 2055 670 3220
rect 950 2055 970 3220
rect 1720 3800 1740 3850
rect 1610 2600 1660 2620
rect 50 1255 100 1275
rect 1525 1255 1575 1275
rect 650 15 670 1180
rect 950 15 970 1180
rect 50 -65 100 -45
rect 1525 -65 1575 -45
<< nsubdiffcont >>
rect 450 5265 500 5285
rect 1125 5265 1175 5285
rect 650 4035 670 5200
rect 950 4035 970 5200
rect 450 3935 500 3955
rect 1125 3935 1175 3955
rect 535 2575 585 2595
rect 1040 2575 1090 2595
rect 645 1345 665 1395
rect 960 1345 980 1395
<< poly >>
rect 1575 5235 1755 5255
rect 0 5220 50 5235
rect 100 5220 150 5235
rect 200 5220 250 5235
rect 300 5220 350 5235
rect 400 5220 450 5235
rect 500 5220 550 5235
rect 735 5220 785 5235
rect 835 5220 885 5235
rect 1075 5220 1125 5235
rect 1175 5220 1225 5235
rect 1275 5220 1325 5235
rect 1375 5220 1425 5235
rect 1475 5220 1525 5235
rect 1575 5220 1625 5235
rect 0 4005 50 4020
rect 100 4005 150 4020
rect 200 4005 250 4020
rect 300 4005 350 4020
rect 400 4005 450 4020
rect 500 4005 550 4020
rect 735 4005 785 4020
rect 835 4005 885 4020
rect 1075 4005 1125 4020
rect 1175 4005 1225 4020
rect 1275 4005 1325 4020
rect 1375 4005 1425 4020
rect 1475 4005 1525 4020
rect 1575 4005 1625 4020
rect 0 3995 1625 4005
rect 0 3990 800 3995
rect 790 3975 800 3990
rect 820 3990 1625 3995
rect 820 3975 830 3990
rect 790 3965 830 3975
rect -45 3910 -5 3920
rect -45 3890 -35 3910
rect -15 3895 -5 3910
rect 155 3910 195 3920
rect 155 3895 165 3910
rect -15 3890 165 3895
rect 185 3895 195 3910
rect 355 3910 395 3920
rect 355 3895 365 3910
rect 185 3890 365 3895
rect 385 3895 395 3910
rect 555 3910 595 3920
rect 555 3895 565 3910
rect 385 3890 450 3895
rect -45 3880 450 3890
rect 0 3865 50 3880
rect 100 3865 150 3880
rect 200 3865 250 3880
rect 300 3865 350 3880
rect 400 3865 450 3880
rect 500 3890 565 3895
rect 585 3890 595 3910
rect 500 3880 595 3890
rect 1030 3910 1070 3920
rect 1030 3890 1040 3910
rect 1060 3895 1070 3910
rect 1230 3910 1270 3920
rect 1230 3895 1240 3910
rect 1060 3890 1125 3895
rect 1030 3880 1125 3890
rect 500 3865 550 3880
rect 1075 3865 1125 3880
rect 1175 3890 1240 3895
rect 1260 3895 1270 3910
rect 1430 3910 1470 3920
rect 1430 3895 1440 3910
rect 1260 3890 1440 3895
rect 1460 3895 1470 3910
rect 1630 3910 1670 3920
rect 1630 3895 1640 3910
rect 1460 3890 1640 3895
rect 1660 3890 1670 3910
rect 1175 3880 1670 3890
rect 1175 3865 1225 3880
rect 1275 3865 1325 3880
rect 1375 3865 1425 3880
rect 1475 3865 1525 3880
rect 1575 3865 1625 3880
rect 735 3240 785 3255
rect 835 3240 885 3255
rect 0 2650 50 2665
rect 100 2650 150 2665
rect 200 2650 250 2665
rect 300 2650 350 2665
rect 400 2650 450 2665
rect 500 2650 550 2665
rect 0 2530 50 2545
rect 100 2530 150 2545
rect 200 2530 250 2545
rect 300 2530 350 2545
rect 400 2530 450 2545
rect 500 2530 550 2545
rect 1075 2650 1125 2665
rect 1175 2650 1225 2665
rect 1275 2650 1325 2665
rect 1375 2650 1425 2665
rect 1475 2650 1525 2665
rect 1575 2650 1625 2665
rect 1075 2530 1125 2545
rect 1175 2530 1225 2545
rect 1275 2530 1325 2545
rect 1375 2530 1425 2545
rect 1475 2530 1525 2545
rect 1575 2530 1625 2545
rect 0 1315 50 1330
rect -45 1305 50 1315
rect -45 1285 -35 1305
rect -15 1300 50 1305
rect 100 1315 150 1330
rect 200 1315 250 1330
rect 300 1315 350 1330
rect 400 1315 450 1330
rect 500 1315 550 1330
rect 100 1305 595 1315
rect 100 1300 165 1305
rect -15 1285 -5 1300
rect -45 1275 -5 1285
rect 155 1285 165 1300
rect 185 1300 365 1305
rect 185 1285 195 1300
rect 155 1275 195 1285
rect 355 1285 365 1300
rect 385 1300 565 1305
rect 385 1285 395 1300
rect 355 1275 395 1285
rect 555 1285 565 1300
rect 585 1285 595 1305
rect 555 1275 595 1285
rect 735 1250 785 2040
rect 835 1250 885 2040
rect 1075 1315 1125 1330
rect 1175 1315 1225 1330
rect 1275 1315 1325 1330
rect 1375 1315 1425 1330
rect 1475 1315 1525 1330
rect 1030 1305 1525 1315
rect 1030 1285 1040 1305
rect 1060 1300 1240 1305
rect 1060 1285 1070 1300
rect 1030 1275 1070 1285
rect 1230 1285 1240 1300
rect 1260 1300 1440 1305
rect 1260 1285 1270 1300
rect 1230 1275 1270 1285
rect 1430 1285 1440 1300
rect 1460 1300 1525 1305
rect 1575 1315 1625 1330
rect 1575 1305 1670 1315
rect 1575 1300 1640 1305
rect 1460 1285 1470 1300
rect 1430 1275 1470 1285
rect 1630 1285 1640 1300
rect 1660 1285 1670 1305
rect 1630 1275 1670 1285
rect 735 1240 885 1250
rect 735 1230 800 1240
rect -130 1220 800 1230
rect 820 1230 885 1240
rect 820 1220 1755 1230
rect -130 1215 1755 1220
rect 0 1200 50 1215
rect 100 1200 150 1215
rect 200 1200 250 1215
rect 300 1200 350 1215
rect 400 1200 450 1215
rect 500 1200 550 1215
rect 735 1210 885 1215
rect 735 1200 785 1210
rect 835 1200 885 1210
rect 1075 1200 1125 1215
rect 1175 1200 1225 1215
rect 1275 1200 1325 1215
rect 1375 1200 1425 1215
rect 1475 1200 1525 1215
rect 1575 1200 1625 1215
rect 0 -15 50 0
rect 100 -15 150 0
rect 200 -15 250 0
rect 300 -15 350 0
rect 400 -15 450 0
rect 500 -15 550 0
rect 735 -15 785 0
rect 835 -15 885 0
rect 1075 -15 1125 0
rect 1175 -15 1225 0
rect 1275 -15 1325 0
rect 1375 -15 1425 0
rect 1475 -15 1525 0
rect 1575 -15 1625 0
<< polycont >>
rect 800 3975 820 3995
rect -35 3890 -15 3910
rect 165 3890 185 3910
rect 365 3890 385 3910
rect 565 3890 585 3910
rect 1040 3890 1060 3910
rect 1240 3890 1260 3910
rect 1440 3890 1460 3910
rect 1640 3890 1660 3910
rect -35 1285 -15 1305
rect 165 1285 185 1305
rect 365 1285 385 1305
rect 565 1285 585 1305
rect 1040 1285 1060 1305
rect 1240 1285 1260 1305
rect 1440 1285 1460 1305
rect 1640 1285 1660 1305
rect 800 1220 820 1240
<< locali >>
rect 440 5285 510 5295
rect 440 5265 450 5285
rect 500 5265 510 5285
rect 440 5255 510 5265
rect -45 5200 -5 5215
rect -45 4035 -35 5200
rect -15 4035 -5 5200
rect -45 3910 -5 4035
rect 55 5200 95 5215
rect 55 4035 65 5200
rect 85 4035 95 5200
rect 55 4025 95 4035
rect 155 5200 195 5215
rect 155 4035 165 5200
rect 185 4035 195 5200
rect 155 4025 195 4035
rect 255 5200 295 5215
rect 255 4035 265 5200
rect 285 4035 295 5200
rect 255 4025 295 4035
rect 355 5200 395 5215
rect 355 4035 365 5200
rect 385 4035 395 5200
rect 355 4025 395 4035
rect 455 5200 495 5255
rect 455 4035 465 5200
rect 485 4035 495 5200
rect 455 3965 495 4035
rect 555 5200 595 5215
rect 555 4035 565 5200
rect 585 4035 595 5200
rect 440 3955 510 3965
rect 440 3935 450 3955
rect 500 3935 510 3955
rect 440 3925 510 3935
rect -45 3890 -35 3910
rect -15 3890 -5 3910
rect -45 3880 -5 3890
rect 155 3910 195 3920
rect 155 3890 165 3910
rect 185 3890 195 3910
rect -125 3850 -5 3860
rect -125 3800 -115 3850
rect -95 3845 -5 3850
rect -95 3820 -35 3845
rect -95 3800 -85 3820
rect -125 3790 -85 3800
rect -45 2680 -35 3820
rect -15 2680 -5 3845
rect -45 2630 -5 2680
rect 55 3845 95 3860
rect 55 2680 65 3845
rect 85 2680 95 3845
rect 55 2650 95 2680
rect 155 3845 195 3890
rect 355 3910 395 3920
rect 355 3890 365 3910
rect 385 3890 395 3910
rect 155 2680 165 3845
rect 185 2680 195 3845
rect 155 2670 195 2680
rect 255 3845 295 3860
rect 255 2680 265 3845
rect 285 2680 295 3845
rect 255 2650 295 2680
rect 355 3845 395 3890
rect 555 3910 595 4035
rect 640 5200 730 5215
rect 640 4035 650 5200
rect 670 4035 700 5200
rect 720 4035 730 5200
rect 640 4025 730 4035
rect 790 5200 830 5215
rect 790 4035 800 5200
rect 820 4035 830 5200
rect 555 3890 565 3910
rect 585 3890 595 3910
rect 355 2680 365 3845
rect 385 2680 395 3845
rect 355 2670 395 2680
rect 455 3845 495 3860
rect 455 2680 465 3845
rect 485 2680 495 3845
rect 455 2650 495 2680
rect 555 3845 595 3890
rect 555 2680 565 3845
rect 585 2680 595 3845
rect 790 3995 830 4035
rect 890 5200 980 5215
rect 890 4035 900 5200
rect 920 4035 950 5200
rect 970 4035 980 5200
rect 890 4025 980 4035
rect 1030 5200 1070 5320
rect 1115 5285 1185 5295
rect 1115 5265 1125 5285
rect 1175 5265 1185 5285
rect 1115 5255 1185 5265
rect 1030 4035 1040 5200
rect 1060 4035 1070 5200
rect 790 3975 800 3995
rect 820 3975 830 3995
rect 555 2670 595 2680
rect 640 3220 730 3235
rect 55 2630 495 2650
rect -45 2620 25 2630
rect -45 2600 -35 2620
rect 15 2600 25 2620
rect -45 2590 25 2600
rect 525 2595 595 2605
rect 525 2575 535 2595
rect 585 2575 595 2595
rect 525 2565 595 2575
rect 55 2545 495 2565
rect -45 2515 -5 2525
rect -45 1350 -35 2515
rect -15 1350 -5 2515
rect -45 1305 -5 1350
rect 55 2515 95 2545
rect 55 1350 65 2515
rect 85 1350 95 2515
rect 55 1335 95 1350
rect 155 2515 195 2525
rect 155 1350 165 2515
rect 185 1350 195 2515
rect -45 1285 -35 1305
rect -15 1285 -5 1305
rect 155 1305 195 1350
rect 255 2515 295 2545
rect 255 1350 265 2515
rect 285 1350 295 2515
rect 255 1335 295 1350
rect 355 2515 395 2525
rect 355 1350 365 2515
rect 385 1350 395 2515
rect 155 1285 165 1305
rect 185 1285 195 1305
rect -45 1260 -5 1285
rect -130 1240 -5 1260
rect 40 1275 110 1285
rect 155 1275 195 1285
rect 355 1305 395 1350
rect 455 2515 495 2545
rect 455 1350 465 2515
rect 485 1350 495 2515
rect 455 1335 495 1350
rect 555 2515 595 2565
rect 555 1350 565 2515
rect 585 1375 595 2515
rect 640 2055 650 3220
rect 670 2055 700 3220
rect 720 2055 730 3220
rect 640 2045 730 2055
rect 790 3220 830 3975
rect 1030 3910 1070 4035
rect 1130 5200 1170 5255
rect 1130 4035 1140 5200
rect 1160 4035 1170 5200
rect 1130 3965 1170 4035
rect 1230 5200 1270 5215
rect 1230 4035 1240 5200
rect 1260 4035 1270 5200
rect 1230 4025 1270 4035
rect 1330 5200 1370 5215
rect 1330 4035 1340 5200
rect 1360 4035 1370 5200
rect 1330 4025 1370 4035
rect 1430 5200 1470 5215
rect 1430 4035 1440 5200
rect 1460 4035 1470 5200
rect 1430 4025 1470 4035
rect 1530 5200 1570 5215
rect 1530 4035 1540 5200
rect 1560 4035 1570 5200
rect 1530 4025 1570 4035
rect 1630 5200 1670 5215
rect 1630 4035 1640 5200
rect 1660 4035 1670 5200
rect 1115 3955 1185 3965
rect 1115 3935 1125 3955
rect 1175 3935 1185 3955
rect 1115 3925 1185 3935
rect 1030 3890 1040 3910
rect 1060 3890 1070 3910
rect 1030 3845 1070 3890
rect 1230 3910 1270 3920
rect 1230 3890 1240 3910
rect 1260 3890 1270 3910
rect 790 2055 800 3220
rect 820 2055 830 3220
rect 790 2045 830 2055
rect 890 3220 980 3235
rect 890 2055 900 3220
rect 920 2055 950 3220
rect 970 2055 980 3220
rect 1030 2680 1040 3845
rect 1060 2680 1070 3845
rect 1030 2670 1070 2680
rect 1130 3845 1170 3860
rect 1130 2680 1140 3845
rect 1160 2680 1170 3845
rect 1130 2650 1170 2680
rect 1230 3845 1270 3890
rect 1430 3910 1470 3920
rect 1430 3890 1440 3910
rect 1460 3890 1470 3910
rect 1230 2680 1240 3845
rect 1260 2680 1270 3845
rect 1230 2670 1270 2680
rect 1330 3845 1370 3860
rect 1330 2680 1340 3845
rect 1360 2680 1370 3845
rect 1330 2650 1370 2680
rect 1430 3845 1470 3890
rect 1630 3910 1670 4035
rect 1630 3890 1640 3910
rect 1660 3890 1670 3910
rect 1630 3880 1670 3890
rect 1430 2680 1440 3845
rect 1460 2680 1470 3845
rect 1430 2670 1470 2680
rect 1530 3845 1570 3860
rect 1530 2680 1540 3845
rect 1560 2680 1570 3845
rect 1530 2650 1570 2680
rect 1130 2630 1570 2650
rect 1630 3850 1750 3860
rect 1630 3845 1720 3850
rect 1630 2680 1640 3845
rect 1660 3820 1720 3845
rect 1660 2680 1670 3820
rect 1710 3800 1720 3820
rect 1740 3800 1750 3850
rect 1710 3790 1750 3800
rect 1630 2630 1670 2680
rect 1600 2620 1670 2630
rect 890 2045 980 2055
rect 1030 2595 1100 2605
rect 1030 2575 1040 2595
rect 1090 2575 1100 2595
rect 1600 2600 1610 2620
rect 1660 2600 1670 2620
rect 1600 2590 1670 2600
rect 1030 2565 1100 2575
rect 1030 2515 1070 2565
rect 635 1395 675 1405
rect 635 1375 645 1395
rect 585 1350 645 1375
rect 555 1345 645 1350
rect 665 1345 675 1395
rect 555 1335 675 1345
rect 950 1395 990 1405
rect 950 1345 960 1395
rect 980 1375 990 1395
rect 1030 1375 1040 2515
rect 980 1350 1040 1375
rect 1060 1350 1070 2515
rect 980 1345 1070 1350
rect 950 1335 1070 1345
rect 1130 2545 1570 2565
rect 1130 2515 1170 2545
rect 1130 1350 1140 2515
rect 1160 1350 1170 2515
rect 1130 1335 1170 1350
rect 1230 2515 1270 2525
rect 1230 1350 1240 2515
rect 1260 1350 1270 2515
rect 355 1285 365 1305
rect 385 1285 395 1305
rect 355 1275 395 1285
rect 555 1305 595 1315
rect 555 1285 565 1305
rect 585 1285 595 1305
rect 40 1255 50 1275
rect 100 1255 110 1275
rect 40 1245 110 1255
rect -45 1185 -5 1240
rect -45 20 -35 1185
rect -15 20 -5 1185
rect -45 5 -5 20
rect 55 1185 95 1245
rect 55 20 65 1185
rect 85 20 95 1185
rect 55 -35 95 20
rect 155 1185 195 1195
rect 155 20 165 1185
rect 185 20 195 1185
rect 155 5 195 20
rect 255 1185 295 1195
rect 255 20 265 1185
rect 285 20 295 1185
rect 255 5 295 20
rect 355 1185 395 1195
rect 355 20 365 1185
rect 385 20 395 1185
rect 355 5 395 20
rect 455 1185 495 1195
rect 455 20 465 1185
rect 485 20 495 1185
rect 455 5 495 20
rect 555 1185 595 1285
rect 1030 1305 1070 1315
rect 1030 1285 1040 1305
rect 1060 1285 1070 1305
rect 790 1240 830 1250
rect 790 1220 800 1240
rect 820 1220 830 1240
rect 555 20 565 1185
rect 585 20 595 1185
rect 555 5 595 20
rect 640 1180 730 1195
rect 640 15 650 1180
rect 670 15 700 1180
rect 720 15 730 1180
rect 640 5 730 15
rect 790 1180 830 1220
rect 790 15 800 1180
rect 820 15 830 1180
rect 40 -45 110 -35
rect 40 -65 50 -45
rect 100 -65 110 -45
rect 40 -75 110 -65
rect 790 -80 830 15
rect 890 1180 980 1195
rect 890 15 900 1180
rect 920 15 950 1180
rect 970 15 980 1180
rect 890 5 980 15
rect 1030 1185 1070 1285
rect 1230 1305 1270 1350
rect 1330 2515 1370 2545
rect 1330 1350 1340 2515
rect 1360 1350 1370 2515
rect 1330 1335 1370 1350
rect 1430 2515 1470 2525
rect 1430 1350 1440 2515
rect 1460 1350 1470 2515
rect 1230 1285 1240 1305
rect 1260 1285 1270 1305
rect 1230 1275 1270 1285
rect 1430 1305 1470 1350
rect 1530 2515 1570 2545
rect 1530 1350 1540 2515
rect 1560 1350 1570 2515
rect 1530 1335 1570 1350
rect 1630 2515 1670 2525
rect 1630 1350 1640 2515
rect 1660 1350 1670 2515
rect 1430 1285 1440 1305
rect 1460 1285 1470 1305
rect 1630 1305 1670 1350
rect 1630 1285 1640 1305
rect 1660 1285 1670 1305
rect 1430 1275 1470 1285
rect 1515 1275 1585 1285
rect 1515 1255 1525 1275
rect 1575 1255 1585 1275
rect 1515 1245 1585 1255
rect 1630 1260 1670 1285
rect 1030 20 1040 1185
rect 1060 20 1070 1185
rect 1030 5 1070 20
rect 1130 1185 1170 1195
rect 1130 20 1140 1185
rect 1160 20 1170 1185
rect 1130 5 1170 20
rect 1230 1185 1270 1195
rect 1230 20 1240 1185
rect 1260 20 1270 1185
rect 1230 5 1270 20
rect 1330 1185 1370 1195
rect 1330 20 1340 1185
rect 1360 20 1370 1185
rect 1330 5 1370 20
rect 1430 1185 1470 1195
rect 1430 20 1440 1185
rect 1460 20 1470 1185
rect 1430 5 1470 20
rect 1530 1185 1570 1245
rect 1530 20 1540 1185
rect 1560 20 1570 1185
rect 1530 -35 1570 20
rect 1630 1240 1755 1260
rect 1630 1185 1670 1240
rect 1630 20 1640 1185
rect 1660 20 1670 1185
rect 1630 5 1670 20
rect 1515 -45 1585 -35
rect 1515 -65 1525 -45
rect 1575 -65 1585 -45
rect 1515 -75 1585 -65
<< viali >>
rect 450 5265 500 5285
rect 450 3935 500 3955
rect -115 3800 -95 3850
rect 650 4035 670 5200
rect 950 4035 970 5200
rect 1125 5265 1175 5285
rect -35 2600 15 2620
rect 535 2575 585 2595
rect 650 2055 670 3220
rect 1125 3935 1175 3955
rect 950 2055 970 3220
rect 1720 3800 1740 3850
rect 1040 2575 1090 2595
rect 1610 2600 1660 2620
rect 645 1345 665 1395
rect 960 1345 980 1395
rect 50 1255 100 1275
rect 650 15 670 1180
rect 50 -65 100 -45
rect 950 15 970 1180
rect 1525 1255 1575 1275
rect 1525 -65 1575 -45
<< metal1 >>
rect -70 5285 1695 5320
rect -70 5265 450 5285
rect 500 5265 1125 5285
rect 1175 5265 1695 5285
rect -70 5200 1695 5265
rect -70 4035 650 5200
rect 670 4035 950 5200
rect 970 4035 1695 5200
rect -70 3955 1695 4035
rect -70 3935 450 3955
rect 500 3935 1125 3955
rect 1175 3935 1695 3955
rect -70 3900 1695 3935
rect -130 3850 210 3865
rect -130 3800 -115 3850
rect -95 3800 210 3850
rect -130 2620 210 3800
rect -130 2600 -35 2620
rect 15 2600 210 2620
rect -130 1275 210 2600
rect 270 3295 1355 3900
rect 270 2595 610 3295
rect 270 2575 535 2595
rect 585 2575 610 2595
rect 270 1430 610 2575
rect 640 3220 980 3255
rect 640 2055 650 3220
rect 670 2055 950 3220
rect 970 2055 980 3220
rect 640 1460 980 2055
rect 1010 2595 1355 3295
rect 1010 2575 1040 2595
rect 1090 2575 1355 2595
rect 270 1395 710 1430
rect 270 1345 645 1395
rect 665 1345 710 1395
rect 270 1310 710 1345
rect 735 1280 885 1460
rect 1010 1430 1355 2575
rect 910 1395 1355 1430
rect 910 1345 960 1395
rect 980 1345 1355 1395
rect 910 1310 1355 1345
rect 1415 3850 1755 3865
rect 1415 3800 1720 3850
rect 1740 3800 1755 3850
rect 1415 2620 1755 3800
rect 1415 2600 1610 2620
rect 1660 2600 1755 2620
rect -130 1255 50 1275
rect 100 1255 210 1275
rect -130 1200 210 1255
rect 635 1200 985 1280
rect 1415 1275 1755 2600
rect 1415 1255 1525 1275
rect 1575 1255 1755 1275
rect 1415 1200 1755 1255
rect -130 1180 1755 1200
rect -130 15 650 1180
rect 670 15 950 1180
rect 970 15 1755 1180
rect -130 -45 1755 15
rect -130 -65 50 -45
rect 100 -65 1525 -45
rect 1575 -65 1755 -45
rect -130 -80 1755 -65
use fcda  fcda_0
timestamp 1697505651
transform 1 0 3236 0 1 -4775
box -224 739 457 9684
<< labels >>
rlabel locali 809 -80 809 -80 5 Ib
rlabel metal1 1050 5320 1050 5320 1 Vcn
rlabel metal1 1755 1250 1755 1250 3 Vcp
rlabel metal1 1755 1220 1755 1220 3 Vbn
rlabel poly 1755 5245 1755 5245 3 Vbp
rlabel metal1 620 -80 620 -80 5 Vn
rlabel metal1 615 5320 615 5320 1 VP
<< end >>
